// What does a hardware wrapper for a module you'd like to test look like?  See below
// for a top-level modeule that serves to send signals to a 7-segment display driver (partically finished).
//
